/***********************************************
 *                                              *
 * Examples for the book Practical UVM          *
 *                                              *
 * Copyright Srivatsa Vasudevan 2010-2016       *
 * All rights reserved                          *
 *                                              *
 * Permission is granted to use this work       * 
 * provided this notice and attached license.txt*
 * are not removed/altered while redistributing *
 * See license.txt for details                  *
 *                                              *
 ************************************************/

`define SLAVE0_MAX  32'hFFFFFFFF
`define SLAVE1_MAX  32'h1FFFFFFF
`define SLAVE2_MAX  32'h2FFFFFFF
`define SLAVE3_MAX  32'h3FFFFFFF
`define SLAVE4_MAX  32'h4FFFFFFF
`define SLAVE5_MAX  32'h5FFFFFFF
`define SLAVE6_MAX  32'h6FFFFFFF
`define SLAVE7_MAX  32'h7FFFFFFF
`define SLAVE8_MAX  32'h8FFFFFFF
`define SLAVE9_MAX  32'h9FFFFFFF
`define SLAVE10_MAX 32'hAFFFFFFF
`define SLAVE11_MAX 32'hBFFFFFFF
`define SLAVE12_MAX 32'hCFFFFFFF
`define SLAVE13_MAX 32'hDFFFFFFF
`define SLAVE14_MAX 32'hEFFFFFFF
`define SLAVE15_MAX 32'hFFFFFF00

`define SLAVE0_MIN  32'h00000000
`define SLAVE1_MIN  32'h10000000
`define SLAVE2_MIN  32'h20000000
`define SLAVE3_MIN  32'h30000000
`define SLAVE4_MIN  32'h40000000
`define SLAVE5_MIN  32'h50000000
`define SLAVE6_MIN  32'h60000000
`define SLAVE7_MIN  32'h70000000
`define SLAVE8_MIN  32'h80000000
`define SLAVE9_MIN  32'h90000000
`define SLAVE10_MIN 32'hA0000000
`define SLAVE11_MIN 32'hB0000000
`define SLAVE12_MIN 32'hC0000000
`define SLAVE13_MIN 32'hD0000000
`define SLAVE14_MIN 32'hE0000000
`define SLAVE15_MIN 32'hF0000000

